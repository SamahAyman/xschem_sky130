**.subckt comparator_multiple
V1 CLK GND PULSE(0 1.8 5n .1n .1n 10n 20n)
V2 A GND PULSE(0 1.8 0 10u 0 0 10u)
V3 B1 GND 0.2
V4 B2 GND 0.4
V5 B3 GND 0.5
V6 B4 GND 0.7
V7 B5 GND 0.9
V8 B6 GND 1
V9 B7 GND 1.1
V10 B8 GND 1.3
V11 B9 GND 1.5
V12 B10 GND 1.7
X1 A B1 CLK Y1 comparator
X2 A B2 CLK Y2 comparator
X3 A B3 CLK Y3 comparator
X4 A B4 CLK Y4 comparator
X5 A B5 CLK Y5 comparator
X6 A B6 CLK Y6 comparator
X7 A B7 CLK Y7 comparator
X8 A B8 CLK Y8 comparator
X9 A B9 CLK Y9 comparator
X10 A B10 CLK Y10 comparator


**** begin user architecture code
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand3/sky130_fd_sc_hd__nand3_1.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfrtp/sky130_fd_sc_hd__dfrtp_1.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor2/sky130_fd_sc_hd__nor2_1.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dlrbn/sky130_fd_sc_hd__dlrbn_1.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a31o/sky130_fd_sc_hd__a31o_2.spice
.include ~/projects/foundry/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_1.spice

**** end user architecture code
**.ends



* expanding   symbol:  /home/ml2/projects/sky130_simulations/comparator.sym # of pins=4
* sym_path: /home/ml2/projects/sky130_simulations/comparator.sym
* sch_path: /home/ml2/projects/sky130_simulations/comparator.sch
.subckt comparator  A B CLK Y
x1 A CLK net3 VGND VNP VPB VPWR net1 sky130_fd_sc_hd__nand3_1
x2 net1 VGND VNP VPB VPWR net2 sky130_fd_sc_hd__inv_1
x3 net2 Y VGND VNP VPB VPWR net5 sky130_fd_sc_hd__nor2_1
x4 net1 CLK B VGND VNP VPB VPWR net3 sky130_fd_sc_hd__nand3_1
x5 A CLK net3 VGND VNP VPB VPWR net1 sky130_fd_sc_hd__nand3_1
x6 net3 VGND VNP VPB VPWR net4 sky130_fd_sc_hd__inv_1
x7 net5 net4 VGND VNP VPB VPWR Y sky130_fd_sc_hd__nor2_1
V1 VGND GND 0
V2 VPWR GND 1.8
V3 VNP GND 0
V4 VPB GND 1.8
.ends

.GLOBAL GND
**** begin user architecture code


.temp 25
vvcc vcc 0 dc 1.8
vvss vss 0 0
.control
tran 5n 10u
plot A CLK Y1+2 Y2+4 Y3+6 Y4+8 Y5+10 Y6+12 Y7+14 Y8+16 Y9+18 Y10+20
.endc


**** end user architecture code
** flattened .save nodes
.end


